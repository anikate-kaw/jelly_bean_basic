package jb_pkg;

  `include "jelly_bean_transaction.sv"
  `include "jelly_bean_seq.sv"
  `include "jb_agent.sv"
  `include "jb_sb.sv"
  `include "jb_env.sv"
  `include "jb_test.sv"

endpackage
